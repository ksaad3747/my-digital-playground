module NOT (
  input  logic a,
  output logic y
);
  assign y = !a;
endmodule : NOT